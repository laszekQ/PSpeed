_ 0 5
system 623937535 18 175 163 3
hollow 1274696703 18 179 152 3
bread 2724009983 24 199 180 3
glass 666129663 20 143 334 3
shield 2786387967 30 241 65 3
