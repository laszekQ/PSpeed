_ 254 6
code 3383652607 18 674 120 10
sword 3678307327 18 378 132 10
browser 1587182079 18 393 15 10
wine 2227890687 18 338 129 10
sword 1945236479 18 199 381 10
mouse 3719501055 18 147 283 10
